module downcounter(
    input rst, c1khz,
    input count, load, 
    input [3:0] pm10,
    input [3:0] pm1,
    input [3:0] ps10,
    input [3:0] ps1,
    output reg [3:0] m10,
    output reg [3:0] m1,
    output reg [3:0] s10,
    output reg [3:0] s1,
    output zero);
    
    // insert your counter code here

endmodule
